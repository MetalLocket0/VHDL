library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;


ENTITY hw4 IS 
   PORT(ipt : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        Z   : OUT STD_LOGIC_VECTOR(6 DOWNTO 0) );
		  
END hw4;


ARCHITECTURE Hdecimal OF hw4 IS
    CONSTANT ZERO : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1000000";  
	 CONSTANT ONE  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1111001";
	 CONSTANT TWO  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100100";
	 CONSTANT THREE: STD_LOGIC_VECTOR(6 DOWNTO 0) := "0110000";
	 CONSTANT FOUR : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0011001";
	 CONSTANT FIVE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0010010";
	 CONSTANT SIX  : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000010";
	 CONSTANT SEVEN: STD_LOGIC_VECTOR(6 DOWNTO 0) := "1111000";
	 CONSTANT EIGHT: STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000000";
	 CONSTANT NINE : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0011000";
	 CONSTANT A    : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001000";
	 CONSTANT B    : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000011";
	 CONSTANT C    : STD_LOGIC_VECTOR(6 DOWNTO 0) := "1000110";
	 CONSTANT D    : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0100001";
	 CONSTANT E    : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0000110";
	 CONSTANT F    : STD_LOGIC_VECTOR(6 DOWNTO 0) := "0001110";
	 CONSTANT BLANK: STD_LOGIC_VECTOR(6 DOWNTO 0) := "1111111";
BEGIN
  const_ipts: PROCESS(ipt)
   BEGIN 
	CASE ipt IS
	WHEN "0000" => Z <= ZERO;
	WHEN "0001" => Z <= ONE;
	WHEN "0010" => Z <= TWO;
	WHEN "0011" => Z <= THREE;
	WHEN "0100" => Z <= FOUR;
	WHEN "0101" => Z <= FIVE;
    WHEN "0110" => Z <= SIX;
	WHEN "0111" => Z <= SEVEN;
	WHEN "1000" => Z <= EIGHT;
	WHEN "1001" => Z <= NINE;
	WHEN "1010" => Z <= A;
	WHEN "1011" => Z <= B;
	WHEN "1100" => Z <= C;
	WHEN "1101" => Z <= D;
	WHEN "1110" => Z <= E;
	WHEN "1111" => Z <= F;
	WHEN OTHERS => Z <= BLANK;
  END CASE;
 END PROCESS;
END Hdecimal;
